module vtml
