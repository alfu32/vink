module vtml

/////////// /////////// import math
/////////// /////////// import term.ui as tui
/////////// /////////// import vxml
/////////// /////////// import arrays
/////////// ///////////
/////////// /////////// [heap]
/////////// /////////// pub struct Event{
/////////// /////////// 	pub mut:
/////////// /////////// 	event_type string
/////////// /////////// 	target     ?&Node
/////////// /////////// }
/////////// ///////////
/////////// /////////// pub fn create(event_type string) Event {
/////////// /////////// 	return Event{
/////////// /////////// 		event_type : event_type
/////////// /////////// 		target: none
/////////// /////////// 	}
/////////// /////////// }
/////////// ///////////
/////////// /////////// pub type EventListener = fn(evt Event)
/////////// ///////////
/////////// /////////// [heap]
/////////// /////////// pub enum StyleKey{
/////////// /////////// 	bg_color
/////////// /////////// 	color
/////////// /////////// 	display
/////////// /////////// 	position
/////////// /////////// 	top
/////////// /////////// 	left
/////////// /////////// 	bottom
/////////// /////////// 	right
/////////// /////////// }
/////////// /////////// pub enum Display{
/////////// /////////// 	inline
/////////// /////////// 	block
/////////// /////////// }
/////////// /////////// pub enum Position{
/////////// /////////// 	absolute
/////////// /////////// 	relative
/////////// /////////// }
/////////// /////////// pub enum LineStyle{
/////////// /////////// 	continuous
/////////// /////////// 	dashed
/////////// /////////// }
/////////// ///////////
/////////// ///////////
/////////// /////////// [heap]
/////////// /////////// pub struct Style{
/////////// /////////// pub mut:
/////////// /////////// 	bg_color u32
/////////// /////////// 	color u32
/////////// /////////// 	display Display
/////////// /////////// 	position Position
/////////// /////////// 	line_style LineStyle
/////////// /////////// 	top ?i32
/////////// /////////// 	left ?i32
/////////// /////////// 	bottom ?i32
/////////// /////////// 	right ?i32
/////////// /////////// 	width ?i32
/////////// /////////// 	height ?i32
/////////// /////////// }
/////////// /////////// pub fn style_default() Style {
/////////// /////////// 	return Style{
/////////// /////////// 		bg_color: 0
/////////// /////////// 		color : 0
/////////// /////////// 		display: .block
/////////// /////////// 		position: .relative
/////////// /////////// 		line_style: .continuous
/////////// /////////// 	}
/////////// /////////// }
/////////// ///////////
/////////// /////////// [heap]
/////////// /////////// struct Node{
/////////// /////////// 	pub mut:
/////////// /////////// 	attributes map[string]string
/////////// /////////// 	children []&Node
/////////// /////////// 	parent_node   ?&Node
/////////// /////////// 	tag_name  string
/////////// /////////// 	listeners map[string][]&EventListener
/////////// /////////// 	style Style
/////////// /////////// 	text string
/////////// /////////// }
/////////// ///////////
/////////// /////////// fn node_create(tag_name string) Node{
/////////// /////////// 	return Node{
/////////// /////////// 		attributes: {}
/////////// /////////// 		children: []
/////////// /////////// 		parent_node: none
/////////// /////////// 		tag_name: tag_name
/////////// /////////// 		listeners: {}
/////////// /////////// 		style: style_default()
/////////// /////////// 		text: ''
/////////// /////////// 	}
/////////// /////////// }
/////////// ///////////
/////////// /////////// fn (this Node) box() Box {
/////////// /////////// 	if this.is_terminal() {
/////////// /////////// 			return Box{
/////////// /////////// 				top : 0
/////////// /////////// 				right: 0
/////////// /////////// 				bottom : 0
/////////// /////////// 				left: this.text.len
/////////// /////////// 			}.pad(1)
/////////// /////////// 	} else {
/////////// /////////// 		return arrays.fold[&Node, Box](this.children,Box{
/////////// /////////// 			top : 0
/////////// /////////// 			right: 0
/////////// /////////// 			bottom : 0
/////////// /////////// 			left: this.text.len
/////////// /////////// 		}.pad(1) , fn(acc Box,n &Node) Box { return acc.add(n.box().pad(1)) } )
/////////// /////////// 	}
/////////// /////////// }
/////////// ///////////
/////////// ///////////
/////////// /////////// fn (this Node) is_terminal() bool {
/////////// /////////// 	return this.children.len == 0
/////////// /////////// }
/////////// /////////// fn (mut this Node) append_child(mut child &Node) {
/////////// /////////// 	if !this.children.contains(child) {
/////////// /////////// 		this.children << child
/////////// /////////// 		child.parent_node = &this
/////////// /////////// 	}
/////////// /////////// }
/////////// ///////////
/////////// /////////// fn (mut this Node) remove_child(mut child &Node) {
/////////// /////////// 	this.children=this.children.filter(it!= child)
/////////// /////////// 	child.parent_node=none
/////////// /////////// }
/////////// ///////////
/////////// /////////// fn (mut this Node) set_attribute(key string,value string) {
/////////// /////////// 	this.attributes[key]=value
/////////// /////////// }
/////////// ///////////
/////////// ///////////
/////////// /////////// fn (this Node) get_attribute(key string) string {
/////////// /////////// 	return this.attributes[key]
/////////// /////////// }
/////////// ///////////
/////////// ///////////
/////////// /////////// fn (mut this Node) remove_event_listener(event_type string,event_listener &EventListener) {
/////////// /////////// 	if !this.listeners.keys().contains(event_type) {
/////////// /////////// 		this.listeners[event_type]=[]
/////////// /////////// 	}
/////////// /////////// 	this.listeners[event_type]=this.listeners[event_type].filter(it!= event_listener)
/////////// /////////// }
/////////// ///////////
/////////// /////////// fn (mut this Node) add_event_listener(event_type string,event_listener &EventListener) {
/////////// /////////// 	if !this.listeners.keys().contains(event_type) {
/////////// /////////// 		this.listeners[event_type]=[]
/////////// /////////// 	}
/////////// /////////// 	this.listeners[event_type] << event_listener
/////////// /////////// }
/////////// ///////////
/////////// /////////// fn (mut this Node) dispatch(event_type string) {
/////////// /////////// 	for listener in this.listeners[event_type] {
/////////// /////////// 		listener(Event{
/////////// /////////// 			target: this
/////////// /////////// 			event_type: event_type
/////////// /////////// 		})
/////////// /////////// 	}
/////////// /////////// }
/////////// /////////// fn (this Node) render(mut ctx &tui.Context,refx i32,refy i32) {
/////////// /////////// 	bx:= this.box()
/////////// /////////// 	ctx.set_bg_color(to_color(this.style.bg_color))
/////////// /////////// 	ctx.set_color(to_color(this.style.color))
/////////// /////////// 	ctx.draw_rect(refx+bx.left,refy+bx.top,refx+bx.right,refy+bx.bottom)
/////////// /////////// 	for child in this.children {
/////////// /////////// 		child.render(mut ctx,refx+bx.left,refy+bx.top)
/////////// /////////// 	}
/////////// /////////// 	ctx.draw_text(refx+bx.left,refy+bx.top,this.text)
/////////// /////////// 	if this.parent_node == none {
/////////// /////////// 		ctx.flush()
/////////// /////////// 	}
/////////// /////////// }
/////////// ///////////
/////////// /////////// pub fn from_vxml_node(vxml_node vxml.Node,parent ?&Node) &Node {
/////////// /////////// 	mut stl:=style_default()
/////////// /////////// 	for attrn,attrv in vxml_node.attributes {
/////////// /////////// 		match attrn {
/////////// /////////// 			"bg_color" { stl.bg_color=attrv.u32() }
/////////// /////////// 			"color" { stl.color=attrv.u32() }
/////////// /////////// 			"display" { stl.display=if attrv=="inline" { Display.inline } else {Display.block} }
/////////// /////////// 			"position" { stl.position=if attrv=="absolute" { Position.absolute } else {Position.relative} }
/////////// /////////// 			"line_style" { stl.line_style=if attrv=="dashed" { LineStyle.dashed } else {LineStyle.continuous} }
/////////// /////////// 			"top" { stl.top=  attrv.u32() }
/////////// /////////// 			"left" { stl.left= attrv.u32() }
/////////// /////////// 			"bottom" { stl.bottom=attrv.u32() }
/////////// /////////// 			"right" { stl.right=attrv.u32() }
/////////// /////////// 			"width" { stl.width=attrv.u32() }
/////////// /////////// 			"height" { stl.height=attrv.u32() }
/////////// /////////// 			else {
/////////// ///////////
/////////// /////////// 			}
/////////// /////////// 		}
/////////// /////////// 	}
/////////// /////////// 	mut vnode := &Node{
/////////// /////////// 		tag_name: vxml_node.name
/////////// /////////// 		parent_node: parent
/////////// /////////// 		attributes: vxml_node.attributes
/////////// /////////// 		style: stl
/////////// /////////// 		text: vxml_node.text
/////////// /////////// 	}
/////////// /////////// 	vnode.children = vxml_node.children.map(from_vxml_node(it,vnode))
/////////// /////////// 	return vnode
/////////// /////////// }
/////////// /////////// pub fn from_xml(xml string) &Node {
/////////// /////////// 	return from_vxml_node(vxml.parse(xml),none)
/////////// /////////// }
